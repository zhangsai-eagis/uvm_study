module tb2;
Data_pkg pkg_1 = new();
  Pkg_a::Data_send_pkg pkg_2;
  initial
      begin
            pkg_2 = new();

          end


endmodule

