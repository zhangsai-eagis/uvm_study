packet m_packet;
  `include m_transation.sv
  `include m_driver.sv
  `include m_env.sv
  `include m_agent.sv
endpacket
